library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;

entity wb_stage is
    port (

        clk                         : in std_logic

    );
end entity;

architecture rtl of wb_stage is

begin


end architecture;