library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity reg_file is
    port (

    );
end entity;

architecture rtl of reg_file is
    signal r0, r1, r2, r3, r4, r5, r6, r7, pc, sp : std_logic_vector(31 downto 0);
begin
    
end architecture;